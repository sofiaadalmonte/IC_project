*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_EX_lpe.spi
#else
.include ../../../work/xsch/JNW_EX.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
*VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
IBP 0 IBPS_5U dc 5u
V0  IBNS_20U 0 dc 1

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save all
.save i(V0) v(IBPS_5U)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1n 10n 1p
write
quit


.endc

.end
